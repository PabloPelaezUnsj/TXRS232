library ieee;
use pablooooooooooooooooo
daleqsovo
