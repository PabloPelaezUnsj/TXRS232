library ieee;
use pablooooooooooooooooo
